`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    12:15:55 03/29/2021 
// Design Name: 
// Module Name:    Registo_de_Flags 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module Registo_de_Flags(
    input clk,
    input [2:0] SEL_F,
    input ESCR_F,
    input [2:0] R_FLAG,
    input bit_maior_peso,
    output S_FLAG
    );


endmodule
